///////////////////////////////////////////////////////////////////////////////
// Module Name: pwm_ramp_adc_subsystem
// 
// Description:
// Implements a PWM ramp-based ADC subsystem with averaging and scaling capabilities.
// The module generates a sawtooth waveform for comparison, captures samples,
// processes them through averaging, and provides multiple output formats.
//
// Inputs:
//   - clk            : System clock
//   - reset          : System reset
//   - compare_match  : Comparator input signal
//   - bin_bcd_select : 2-bit output format selector
//
// Outputs:
//   - pwm_out       : PWM output signal
//   - adc_outputs   : 16-bit processed ADC output
//
// Internal Signals:
//   - u8_raw_data    : 8-bit raw ADC sample
//   - ave_data       : 16-bit averaged data
//   - scaled_ave_hex : Scaled averaged data in hex
//   - scaled_ave_dec : Scaled averaged data in BCD
//   - ready_pulse    : Sample capture trigger
//
// Operation:
//   1. Sawtooth generator produces 100Hz reference waveform
//   2. Sample capture triggers on comparator transitions
//   3. Raw samples are averaged over 64 samples (2^6)
//   4. Averaged data is scaled by factor of 120 with +150 offset
//   5. Output format selected via bin_bcd_select:
//      00: Scaled average (hex)
//      01: Scaled average (BCD)
//      10: Raw ADC data
//      11: Averaged data
//
// Note: Averager configured for 6-bit power (64 samples) to improve resolution
//       while maintaining reasonable response time
///////////////////////////////////////////////////////////////////////////////


module pwm_ramp_adc_subsystem(
    input logic clk,
    input logic reset,
    input logic compare_match,
    input logic [1:0] bin_bcd_select, 

    output logic   pwm_out,
    output logic [15:0] adc_outputs
);
    
            
    logic [7:0] u8_raw_data;              // Raw ADC data
    logic [15:0] ave_data;
    logic [15:0] scaled_data;
    logic [15:0] scaled_ave_hex; // Scaled ADC data for display, plus pipelinging register
    logic [15:0] scaled_ave_dec; // Scaled ADC data for display, plus pipelinging register

    // Output assignments
    assign raw_adc_data_out = u8_raw_data;
    assign ave_adc_data_out = ave_data;
    assign scaled_adc_data_out = scaled_data;



    logic pwm_out_internal;
    logic [7:0] R2R_out_internal;
    
    logic sawtooth_en;
    assign sawtooth_en = 1;
    // Instantiate the triangle_generator module
    sawtooth_waveform #(
        .WIDTH(8),           // Bit width for duty_cycle (e.g. 8)
        .CLOCK_FREQ(100_000_000), // System clock frequency in Hz (e.g. 100_000_000)
        .WAVE_FREQ(100.0)    // Desired triangle wave frequency in Hz (e.g. 1.0)
    ) sawtooth_pwm_inst (
        .clk(clk),           // Connect to system clock
        .reset(reset),       // Connect to system reset
        .enable(sawtooth_en), // Connect to enable signal
        .pwm_out(pwm_out_internal), // Connect to PWM output signal
        .R2R_out(R2R_out_internal)  // Connect to R2R ladder header, can leave empty if 
    );  
    
    assign pwm_out = pwm_out_internal;
    
    // added sample_capture generated by Claude ai
    // falling edge detector included no need for inverter
    
    logic ready_pulse;
    sample_capture SAMPLE_CAPTURE
    (
        .clk(clk),
        .reset(reset),
        .compare_match(compare_match),
        .R2R_input(R2R_out_internal),
        .u8_raw_data(u8_raw_data),
        .ready_pulse(ready_pulse)
        
    );
    
    
    // average data is scaled and stored
    always_ff @(posedge clk) begin
        if (reset)
            scaled_ave_hex <= '0;
        else if (ready_pulse)
            scaled_ave_hex <= (ave_data * 120 + 150);  // Approximate scaling factor
    end
    
    bin_to_bcd  DECIMAL_CONVERTER
    (
        .clk(clk),
        .reset(reset),
        .bin_in(scaled_ave_hex),
        .bcd_out(scaled_ave_dec)
    );


        
    // average
    averager #(
        .power(6), // 2**(power) samples, default is 2**8 = 256 samples (4^4 = 256 samples, adds 4 bits of ADC resolution)
        .N(12)     // # of bits to take the average of
    ) AVERAGER (
        .reset(reset),
        .clk(clk),
        .EN(ready_pulse),
        .Din(u8_raw_data),
        .Q(ave_data)
    );
    
 
 logic [15:0] adc_mux_outputs;

 always_comb begin
    case(bin_bcd_select)
        2'b00: adc_mux_outputs= scaled_ave_hex;  // averaged ADC with extra 4 bits
        2'b01: adc_mux_outputs = scaled_ave_dec;  // averaged and scaled voltage
        2'b10: adc_mux_outputs = u8_raw_data;  // raw ADC (12-bits)
        2'b11: adc_mux_outputs = ave_data;
        default: adc_mux_outputs = scaled_ave_hex;  // Default case: output all zeros
    endcase
  end
  
  assign  adc_outputs = adc_mux_outputs;   
  
endmodule
      